module display_matrix(clk, rst, pattern_id, dot_row, dot_col);
	input				clk, rst;
	input		[3:0]	pattern_id;
	output reg	[7:0]	dot_row, dot_col;
	reg			[2:0]	row_cnt;

	always @(posedge clk or negedge rst) begin
		if (!rst) begin
			dot_row <= 0;
			dot_col <= 0;
			row_cnt <= 0;
		end
		else begin
			case ({row_cnt, pattern_id})
				7'b000_0001: dot_col <= 8'b00000000;
				7'b001_0001: dot_col <= 8'b00000000;
				7'b010_0001: dot_col <= 8'b00000000;
				7'b011_0001: dot_col <= 8'b00000000;
				7'b100_0001: dot_col <= 8'b00010000;
				7'b101_0001: dot_col <= 8'b00000000;
				7'b110_0001: dot_col <= 8'b00000000;
				7'b111_0001: dot_col <= 8'b00000000;

				7'b000_0010: dot_col <= 8'b00000000;
				7'b001_0010: dot_col <= 8'b00000000;
				7'b010_0010: dot_col <= 8'b00000000;
				7'b011_0010: dot_col <= 8'b00011000;
				7'b100_0010: dot_col <= 8'b00011000;
				7'b101_0010: dot_col <= 8'b00000000;
				7'b110_0010: dot_col <= 8'b00000000;
				7'b111_0010: dot_col <= 8'b00000000;

				7'b000_0011: dot_col <= 8'b00000000;
				7'b001_0011: dot_col <= 8'b00000000;
				7'b010_0011: dot_col <= 8'b00000000;
				7'b011_0011: dot_col <= 8'b00110000;
				7'b100_0011: dot_col <= 8'b00101000;
				7'b101_0011: dot_col <= 8'b00010000;
				7'b110_0011: dot_col <= 8'b00000000;
				7'b111_0011: dot_col <= 8'b00000000;

				7'b000_0100: dot_col <= 8'b00000000;
				7'b001_0100: dot_col <= 8'b00000000;
				7'b010_0100: dot_col <= 8'b00000000;
				7'b011_0100: dot_col <= 8'b00010000;
				7'b100_0100: dot_col <= 8'b00101000;
				7'b101_0100: dot_col <= 8'b00010000;
				7'b110_0100: dot_col <= 8'b00000000;
				7'b111_0100: dot_col <= 8'b00000000;

				7'b000_0101: dot_col <= 8'b00000000;
				7'b001_0101: dot_col <= 8'b00000000;
				7'b010_0101: dot_col <= 8'b00000000;
				7'b011_0101: dot_col <= 8'b00011000;
				7'b100_0101: dot_col <= 8'b00100100;
				7'b101_0101: dot_col <= 8'b00011000;
				7'b110_0101: dot_col <= 8'b00000000;
				7'b111_0101: dot_col <= 8'b00000000;

				7'b000_0110: dot_col <= 8'b00000000;
				7'b001_0110: dot_col <= 8'b00000000;
				7'b010_0110: dot_col <= 8'b00011000;
				7'b011_0110: dot_col <= 8'b00100100;
				7'b100_0110: dot_col <= 8'b00010100;
				7'b101_0110: dot_col <= 8'b00001000;
				7'b110_0110: dot_col <= 8'b00000000;
				7'b111_0110: dot_col <= 8'b00000000;

				7'b000_0111: dot_col <= 8'b00000000;
				7'b001_0111: dot_col <= 8'b00000000;
				7'b010_0111: dot_col <= 8'b00000000;
				7'b011_0111: dot_col <= 8'b00000000;
				7'b100_0111: dot_col <= 8'b00111000;
				7'b101_0111: dot_col <= 8'b00000000;
				7'b110_0111: dot_col <= 8'b00000000;
				7'b111_0111: dot_col <= 8'b00000000;

				7'b000_1000: dot_col <= 8'b00000000;
				7'b001_1000: dot_col <= 8'b00000000;
				7'b010_1000: dot_col <= 8'b00110000;
				7'b011_1000: dot_col <= 8'b00110000;
				7'b100_1000: dot_col <= 8'b00001100;
				7'b101_1000: dot_col <= 8'b00001100;
				7'b110_1000: dot_col <= 8'b00000000;
				7'b111_1000: dot_col <= 8'b00000000;

				7'b000_1001: dot_col <= 8'b00000000;
				7'b001_1001: dot_col <= 8'b00000000;
				7'b010_1001: dot_col <= 8'b00000000;
				7'b011_1001: dot_col <= 8'b00010000;
				7'b100_1001: dot_col <= 8'b00001000;
				7'b101_1001: dot_col <= 8'b00111000;
				7'b110_1001: dot_col <= 8'b00000000;
				7'b111_1001: dot_col <= 8'b00000000;

				7'b000_1010: dot_col <= 8'b00000000;
				7'b001_1010: dot_col <= 8'b00000000;
				7'b010_1010: dot_col <= 8'b01001000;
				7'b011_1010: dot_col <= 8'b00000100;
				7'b100_1010: dot_col <= 8'b01000100;
				7'b101_1010: dot_col <= 8'b00111100;
				7'b110_1010: dot_col <= 8'b00000000;
				7'b111_1010: dot_col <= 8'b00000000;

				7'b000_1011: dot_col <= 8'b00000000;
				7'b001_1011: dot_col <= 8'b00000000;
				7'b010_1011: dot_col <= 8'b00010000;
				7'b011_1011: dot_col <= 8'b01000100;
				7'b100_1011: dot_col <= 8'b00000010;
				7'b101_1011: dot_col <= 8'b01000010;
				7'b110_1011: dot_col <= 8'b00111110;
				7'b111_1011: dot_col <= 8'b00000000;

				7'b000_1100: dot_col <= 8'b00000000;
				7'b001_1100: dot_col <= 8'b00000000;
				7'b010_1100: dot_col <= 8'b00101000;
				7'b011_1100: dot_col <= 8'b01000000;
				7'b100_1100: dot_col <= 8'b00100100;
				7'b101_1100: dot_col <= 8'b00001110;
				7'b110_1100: dot_col <= 8'b00000000;
				7'b111_1100: dot_col <= 8'b00000000;

				7'b000_1101: dot_col <= 8'b00000000;
				7'b001_1101: dot_col <= 8'b00000000;
				7'b010_1101: dot_col <= 8'b00111000;
				7'b011_1101: dot_col <= 8'b00000000;
				7'b100_1101: dot_col <= 8'b00010000;
				7'b101_1101: dot_col <= 8'b00010000;
				7'b110_1101: dot_col <= 8'b00010000;
				7'b111_1101: dot_col <= 8'b00000000;

				7'b000_1110: dot_col <= 8'b00000000;
				7'b001_1110: dot_col <= 8'b00000000;
				7'b010_1110: dot_col <= 8'b00000000;
				7'b011_1110: dot_col <= 8'b00110100;
				7'b100_1110: dot_col <= 8'b00100100;
				7'b101_1110: dot_col <= 8'b00101100;
				7'b110_1110: dot_col <= 8'b00000000;
				7'b111_1110: dot_col <= 8'b00000000;

				7'b000_1111: dot_col <= 8'b00000000;
				7'b001_1111: dot_col <= 8'b00000000;
				7'b010_1111: dot_col <= 8'b00000000;
				7'b011_1111: dot_col <= 8'b01000000;
				7'b100_1111: dot_col <= 8'b00010000;
				7'b101_1111: dot_col <= 8'b11001110;
				7'b110_1111: dot_col <= 8'b00000000;
				7'b111_1111: dot_col <= 8'b00000000;

				default: dot_col <= 0;
			endcase
			case (row_cnt)
				3'd0: dot_row <= 8'b01111111;	
				3'd1: dot_row <= 8'b10111111;	
				3'd2: dot_row <= 8'b11011111;	
				3'd3: dot_row <= 8'b11101111;	
				3'd4: dot_row <= 8'b11110111;	
				3'd5: dot_row <= 8'b11111011;	
				3'd6: dot_row <= 8'b11111101;	
				3'd7: dot_row <= 8'b11111110;	
			endcase
			row_cnt <= row_cnt + 1;
		end
	end
endmodule
